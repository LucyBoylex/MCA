BZh91AY&SY��B A�_�Ryg���g������`���y}2�� �y����f��8 �al-� DJ��`�on�'�iZ�e���h	�&��$����S�i�6�i�=OPdh)T��h� 1� ɐ�j��%H        )�EU20 F   &# D��z	�T�M��`C�4�����A )@& f�������4bmw"��;���s��H����T�(l�;���TR�iB�~�]���������۫l4�JS[EO|K�QHYE�p�u� ���L��l�,"g�� M6�c�^z��Y��V'��T$8w�8���7j���s��w�W�j�AJ����$�����me@M��� M�2�b�We'l�^�p�f�D����@�	H�n6um��pD��n�hm�/1ݤ��pJT�G#Vu+7dSe��gkQ<�kH��2���!�j��r�M<����ْ�-�Z:�֍oET �)<���۪�T����c1U�˞;�gX�F�W[�d�����FըIVHa���9�T� �+���Ww�)JJ΅D��R]T�Υ��n�+�K�kv�7 �g��5ܳ{��a��x*\���3J1a.����H�/$��5��ͩ+��l��QK�1�Ҧ��L�I�[f$Lt�A2����$��P%q�1b�0:��2����h�f�L��c��2�i��u�q"ִҥ�e��f�V]uX��{�<^\����$��{R�D,ju�#�:�K�����iP\s����t2C ��	q3�h��	�#m������k� I"�@t[D��(�H���L\�"Gl�pt�8�`aqQc�,e��
�h+&M�Vb�ѭkEPUh���km�AB���ٙ҂n,Ub��6B#Z������*D�UuP�]A	 �ا��b2� b%"-�TF�m�K�r���i%���t�aa`P�B�ITj:rX�3&zdӲub��IX���Z�s��;l拴��]cad���s}*���V�Upm�!�S{i�'������WǛ�
�O�T6\���՝4�ν�xNl�<;�-A�u5x'�>5S}�6(�T6C��Y&EV�}�V�ͬ����}�K�ʧY�%���ʐ�3�S���7�����Tw�ފ�r��ݳ�f���)��li9=:��<��Ǒ}�glVVN�2Ul�k�ͬ�Yt���8&B��WʗS%UU�]ƕ�n�Wݻ6+d��ԩ��_
ʻ�F��s;Z�٭U�r2��yDN��-�gefTܻ�ܻ�ζ:�۰�n����5v��\y�V6�T&���Z����J����S��H�$�����@I�l�I!h8�]o~7�Qg�F�@�����>(�E F�����ߎ#�(�����B��B�DF"�DEF�U�d�-���j'͗��(�T@�wdcr��3��*�El�IR���ٗr�/��.�\.���u�ASC� ��x�1�_������]���u�p)�m9��"��Q�a�٠���h�K(n���7%Cl�������lѰ����gB�����C���j�)�܇v�����adR@��4�h�Z��o����P+QU�d1x��L�B:�i���E	b(�P8dp���&b��R��Z�{9��.���!���*���:�`$�U���Ie1a��D�PI�%1�B��Rj�\k�|�����Ʉ��Y�K���L[Y�clXKm�����6G��ӔO4,�a�����*	c�!�Ѕs�U)*��I��-\X�co�5�tj}i��,�y��;�%�ߜ6$A"���<�in۹&L�����l���J�d�qE��n��rp��.���,W���U�z�:lC�|c�8�JZ��yt��B��<Z��'Bh<i��M���-�,�Cͅ��u$��gN��V���J
|M�K�A���o�l�P��8ӣ!GE�VE$�-�=k#�.Ƣ�S^�Yx����.���c�B0H���R�%II�U��u]mK��ç2慮���&9a�,4E�	����̂	@�!,��2  RPc��84.��U4���;�ZK��~k~��{İ�0�x8x���fܰ|R=31�e�T@�d8��
3���J�����'B�b����P+FE)��Aa����9za�փ��I
�̣q��_IĴ9��x���Pj��[+;��"#MidiV�UPQD=�
;�
S����Vp=��2*��2Yl�DdI#icum�ۗ+���6HohўzŌ��oua�U���]@�S��z�1f�m-�ٱ`#��9GGR�DU�Hy<�����8W��:�<d0ϋu�v�0(��4�G�T��!�F�� 4�YG ��KM������L��>2&�.�:4k�Mgn<�������B�0�}!�z^D�vl���T�w$�(���v��V9Kf�z@se;�V@9��Q	 ��r��e4-2��Q��4�M�U�U�h�nQr�@:j�vx�~f6eʹW"K�Ŷ
���7�s2�I�����u�3&�QOC�-,/L��nYFb�q @���Gr���R��u,C�$�(�Q��s�7Z|=$�Y}���n��0���4!����i�i.��g=�
	VeJ6+��
���7���az�2H�����a�1�О�23@���9
�Y��Yg��͇ٗM `����T��n�e�](8�Bk��4C��ee{�74�8o�N�;�`��\��e�p�窬��ve�!�Vw}-y�-�j�}����Kx��HhE���vIDi�BFT)F�ZAh�EQj�j�u��܀�Hԕ�%W��C˖��A��I7x�V%���m��߃�^H��Çg]i�B����Ôml�f�z�e� iѣ!�8ٝhσ�3UU%S��!���Xx/�����(�mօ�g��\�w�s��,<LV��G<M��q��i�����Kf��*a ׾�5uÕu��������u��I9,Z9��
U���e��˄dH--���
R�2Q��� i��m:� {�qfz����}rK4h�i�S�@�:%�8��p3�.Kq�N��D�a��P��ޛ�	N,7�4�-S�^�ڏ@2�d��!�e�μ�2�7��� �6x�g(��A����eN���f;:p��pg�HH�HFH�$R!��DL�Isv�(TG�����R�U�xˊJGWr6�d�d�_;�@3�r�w.U�(��d�����(~;ԙrdє�c�PzNTfwq&d̑�:j�tU�!�T>H���+5F���^p��-tY��#B�I�5I#w"@��N7�6Ï|��ⷺ�.��V�e������8��\��ʙ^#B�l1C��:ȕ�K:��C�����C�w�gM�]C{�ݪ�^c2c<=5��n�Ȋ�ke��
+�r��x"�0�#"�(H�!s*@R%�B�))���Q�Y�ա���욕]\���L�q-�t�Q�&^��d�#�0�0J�jw����S
B�H��&�|���FX��=%tK<���k�C}�l�	��4a-�x�ͼ��/^���ɇI�$����v9 i���y��C�ְV['9<��d<l��ˣ@�ƃG`+��<9[Y���2Y���ɉR4lbx�w���nrF䑌�T��7.K ܙ1-S$i��$���gΓ�$�. 8��ɰ��A�s�x�r
ٌ��Bd�����tqb+�S9}^$�N�NL����.N�VC��=/o1l��Q�1��f�$��a�e�l��L�h"T'52�@�N�(Z)�.�Y��=&�B�$�I ETR�O:*)���G�b�t�����J͢��Q�>2Cc@�#Q�"U4
�+Q4f�`�b�@ +�j��)��� ����H�XERb�`�X�� ,6@�c ��"*� YdR�# � � ��B� Z �2*H#���Ѣ1G&j�@��F���d�p;Y��>	� ��*ȳ+nu����������ew+�7����)=߶�o��~�T��xon�06���������v;Y��:�@��!��q��K�՗+�BHH��x�Y.���^�X��QM�QO�)Jha�u�M�o�w�'�6's�����p:�!�7:���J*)����Kτ8�̿I��H6\C�S��P�<!�J��a�sg|j��99MJQ�%`S8!$$t������a��]3�p3s�EAN0E0�@� ,"1&�%X�0�d��$���	"�b��"�F �,�1D� �#�[!��>X��D�lq6"���"��+�l9�'a0������l&X�BQR��a%0�
�h�v�Ό��|n�l|���q�=�_����g
(���R�&���,,H������U��IG��p��5�z�[���g٥MȨ����� 
��L���^LLג�f���`�(7w��-ױ�ރ�N���9Qh`��ĸ�p��{T*�v�%�g(���m	Vى[*Z
*B�\�)b�i΅0��J%@S����S.������b�B��G�9	���xZ*)�}+�[���B3�NF�訧����ӱdG���|�y��7"������h�&��C� x����4����QJӈ�r��!���( q<�2*)��c$�QH�7� ��:��жfq2(q"�꼐�x��
b-�pX���QYeU�Rf!���/�}�I	1���rw|��-��4	W)�䩠Wr.d$��m�-�8�V3��k��&�������E.>�HZCv��.�>aTRp��Ǝ@�`*�o7:�NdTR�ٸ�8Y#-�Tn�O�>��H�Y�����j���rE8P���B